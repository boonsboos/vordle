module main

import game

fn main() {
	println("welcome to vordle.")
	game.game()
}